
class sample;
  	rand unsigned int data;
  	int q[$];
  function pre_randomize();
    if(q.size()==8)
      q.delete();
  endfunction
  function post_randomize();
    q.pushback(a);
  endfunction
endclass
module top;
  sample s=new();
  initial begin
    repeat(5);
    assert(s.randomize());
  end
endmodule
=====================================RESULT=================================
Data=3, Q='{3} 
Data=22, Q='{3, 22} 
Data=1, Q='{3, 22, 1} 
Data=9, Q='{3, 22, 1, 9} 
Data=13, Q='{3, 22, 1, 9, 13} 
Data=7, Q='{3, 22, 1, 9, 13, 7} 
Data=16, Q='{3, 22, 1, 9, 13, 7, 16} 
Data=18, Q='{3, 22, 1, 9, 13, 7, 16, 18} 
Data=29, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29} 
Data=26, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26} 
Data=15, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15} 
Data=31, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31} 
Data=31, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31} 
Data=30, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30} 
Data=26, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30} 
Data=27, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27} 
Data=20, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20} 
Data=3, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20} 
Data=8, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8} 
Data=6, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6} 
Data=0, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0} 
Data=17, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=8, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=29, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=13, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=31, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=15, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=1, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17} 
Data=25, Q='{3, 22, 1, 9, 13, 7, 16, 18, 29, 26, 15, 31, 30, 27, 20, 8, 6, 0, 17, 25} 
Data=8, Q='{8} 
Data=30, Q='{8, 30} 
Data=23, Q='{8, 30, 23} 
Data=14, Q='{8, 30, 23, 14} 
Data=9, Q='{8, 30, 23, 14, 9} 
Data=23, Q='{8, 30, 23, 14, 9} 
Data=24, Q='{8, 30, 23, 14, 9, 24} 
Data=30, Q='{8, 30, 23, 14, 9, 24} 
Data=30, Q='{8, 30, 23, 14, 9, 24} 
Data=22, Q='{8, 30, 23, 14, 9, 24, 22} 
Data=19, Q='{8, 30, 23, 14, 9, 24, 22, 19} 
Data=15, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15} 
Data=13, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13} 
Data=25, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25} 
Data=29, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29} 
Data=31, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29, 31} 
Data=22, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29, 31} 
Data=10, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29, 31, 10} 
Data=31, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29, 31, 10} 
Data=30, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29, 31, 10} 
Data=26, Q='{8, 30, 23, 14, 9, 24, 22, 19, 15, 13, 25, 29, 31, 10, 26} 
